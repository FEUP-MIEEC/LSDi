library verilog;
use verilog.vl_types.all;
entity adder4b_tb is
end adder4b_tb;
