library verilog;
use verilog.vl_types.all;
entity lsdalu_testbench is
end lsdalu_testbench;
