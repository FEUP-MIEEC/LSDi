library verilog;
use verilog.vl_types.all;
entity NOR8_MXILINX_detFlags is
    port(
        I0              : in     vl_logic;
        I1              : in     vl_logic;
        I2              : in     vl_logic;
        I3              : in     vl_logic;
        I4              : in     vl_logic;
        I5              : in     vl_logic;
        I6              : in     vl_logic;
        I7              : in     vl_logic;
        O               : out    vl_logic
    );
end NOR8_MXILINX_detFlags;
