library verilog;
use verilog.vl_types.all;
entity addsub4b_tb is
end addsub4b_tb;
