library verilog;
use verilog.vl_types.all;
entity fulladder_tb is
end fulladder_tb;
